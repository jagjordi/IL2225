../SOURCE/tb_FIR.vhd